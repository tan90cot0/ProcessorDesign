LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;
    USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PRGM_TB IS 

END ENTITY;

ARCHITECTURE BEV OF PRGM_TB IS

SIGNAL ADDRESS : STD_LOGIC_VECTOR(5 DOWNTO 0):="000000";
SIGNAL DATAOUT : STD_LOGIC_VECTOR(31 DOWNTO 0);

COMPONENT PRGM IS
    PORT(
         ADDRESS : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
         DATAOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
         );
END COMPONENT;

BEGIN

  UUT: PRGM PORT MAP(ADDRESS, DATAOUT);

  PROCESS
  BEGIN
    ADDRESS<="111111";
    WAIT FOR 100 ns;
    ADDRESS<="111110";
    WAIT FOR 100 ns;
    ADDRESS<="111101";
    WAIT FOR 100 ns;
    ADDRESS<="111100";
    WAIT FOR 100 ns;
    ADDRESS<="000011";
    WAIT FOR 100 ns;
    ADDRESS<="000100";
    WAIT FOR 100 ns;
    ADDRESS<="000101";
    WAIT FOR 100 ns;
    
    ASSERT FALSE REPORT "Test done. Open EPWave to see signals." SEVERITY NOTE;
    WAIT;
  END PROCESS;

END BEV;
