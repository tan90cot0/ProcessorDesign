LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;
    USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PRGM IS
  PORT(
       ADDRESS : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
       DATAOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
       );
END ENTITY;

ARCHITECTURE BEV OF PRGM IS

TYPE MEM IS ARRAY (63 DOWNTO 0) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL MEMORY : MEM := (x"00000010",x"00000011",x"00000000", x"00000100",others => x"00000000");
SIGNAL ADDR : INTEGER RANGE 0 TO 63;

BEGIN
    ADDR<=CONV_INTEGER(ADDRESS);
    DATAOUT<=MEMORY(ADDR);
END BEV;